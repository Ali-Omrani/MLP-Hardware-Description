----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:36:09 12/15/2017 
-- Design Name: 
-- Module Name:    ROM - n1_1 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
use work.fixed_point_package.all;
package fixed_point_array_pkg is
	type fixed_point_array is array(natural range <>) of fixed_point;
end package;

library ieee;
use ieee.std_logic_1164.all;
use work.fixed_point_array_pkg.all;
use work.fixed_point_package.all;

entity ROM is
	generic(
		address_size : integer;
		entry_length : integer
	);
	port(
		clk	: in std_logic;
		en 	: in std_logic;
		address : in integer;
		ROM_data	: out fixed_point_array (0 to address_size-1)
	);
end ROM;

architecture weight_L1 of ROM is

	type rom_type is array (0 to address_size-1) of fixed_point_array (0 to entry_length-1);
	signal rom : rom_type:=(
(('0', "000000000000110"),('0', "000000000001010"),('1', "000000000011010"),('0', "000000000000111"),('0', "000000001000111"),('1', "000000000100101"),('0', "000000000010111"),('1', "000000000000011"),('0', "000000001100100"),('0', "000000000001100"),('0', "000000000010000"),('0', "000000000110001"),('0', "000000000101110"),('1', "000000001000010"),('0', "000000001011010"),('0', "000000000000010"),('1', "000000000010110"),('0', "000000000000110"),('0', "000000000001010"),('1', "000000010100000"),('1', "000000010101010"),('1', "000000010011011"),('1', "000000000001001"),('0', "000000000000001"),('0', "000000000111101"),('0', "000000000111100"),('1', "000000000100000"),('1', "000000000110111"),('1', "000000000100111"),('1', "000000011011010"),('0', "000000000101110"),('0', "000000000111100"),('0', "000000000100100"),('1', "000000000010011"),('1', "000000001111010"),('0', "000000000001010"),('0', "000000011001100"),('1', "000000001101010"),('1', "000000000001100"),('1', "000000001011101"),('1', "000000000110001"),('1', "000000000011101"),('0', "000000001111010"),('1', "000000001111000"),('1', "000000000010100"),('1', "000000010000001"),('1', "000000001110000"),('0', "000000001010011"),('0', "000000000110000"),('1', "000000001000101"),('0', "000000000011101"),('0', "000000001000100"),('0', "000000000010110"),('1', "000000000001000"),('0', "000000000001110"),('0', "000000000011011"),('0', "000000001101010"),('0', "000000000001111"),('0', "000000000111000"),('1', "000000001011101"),('0', "000000000110001"),('0', "000000000011100"),('1', "000000011010001")),
 ------------------------------- 
(('0', "000000001011011"),('1', "000000001100010"),('0', "000000000111011"),('1', "000000000100011"),('0', "000000001010110"),('0', "000000000110100"),('0', "000000001011111"),('0', "000000001101011"),('1', "000000010001111"),('1', "000000001010011"),('0', "000000000110100"),('1', "000000000101011"),('0', "000000010000111"),('0', "000000000110000"),('1', "000000001001101"),('0', "000000001011011"),('0', "000000000100110"),('1', "000000010001000"),('0', "000000001010100"),('1', "000000000100000"),('0', "000000001111111"),('1', "000000000110100"),('1', "000000001100101"),('0', "000000010001001"),('1', "000000001010110"),('0', "000000000000101"),('1', "000000001100010"),('1', "000000000101000"),('0', "000000001110010"),('0', "000000000000011"),('1', "000000011010010"),('1', "000000000000110"),('0', "000000000100111"),('1', "000000100100011"),('0', "000000000101110"),('1', "000000000101110"),('1', "000000011001111"),('0', "000000010101001"),('1', "000000100010001"),('0', "000000000000100"),('1', "000000001110101"),('1', "000000010010011"),('0', "000000001010100"),('0', "000000010000010"),('0', "000000010111000"),('0', "000000100001111"),('0', "000000001110101"),('0', "000000001110100"),('0', "000000100000111"),('1', "000000000101101"),('0', "000000000101100"),('0', "000000100000000"),('1', "000000000001010"),('0', "000000000000101"),('0', "000000000001001"),('0', "000000010100010"),('0', "000000001100000"),('1', "000000100000100"),('1', "000000001011101"),('0', "000000000010001"),('1', "000000010010011"),('1', "000000001001011"),('0', "000000000000111")),
 ------------------------------- 
(('1', "000000000011111"),('1', "000000000000011"),('1', "000000010100011"),('1', "000000000100110"),('0', "000000001001110"),('0', "000000000001110"),('1', "000000001000000"),('1', "000000001111111"),('1', "000000000100100"),('1', "000000000110000"),('0', "000000001111010"),('1', "000000000001000"),('0', "000000001010100"),('1', "000000010000000"),('1', "000000011111011"),('0', "000000001000101"),('0', "000000000000100"),('1', "000000010001100"),('0', "000000010011001"),('0', "000000000001111"),('1', "000000001100101"),('1', "000000000111101"),('1', "000000001010101"),('1', "000000001001000"),('0', "000000000111010"),('1', "000000000101101"),('0', "000000000111001"),('1', "000000000111000"),('0', "000000001110100"),('0', "000000000111010"),('0', "000000001001111"),('1', "000000000110001"),('0', "000000000100100"),('1', "000000000010011"),('0', "000000000001001"),('1', "000000011000110"),('1', "000000010100110"),('0', "000000001010001"),('0', "000000010000100"),('0', "000000000111100"),('0', "000000001111101"),('0', "000000000101101"),('0', "000000011101100"),('0', "000000011101001"),('0', "000000000011111"),('0', "000000000111000"),('1', "000000001101011"),('0', "000000010001111"),('1', "000000001100111"),('1', "000000001100000"),('0', "000000001100101"),('0', "000000000000101"),('0', "000000001001101"),('0', "000000000001101"),('0', "000000010000101"),('1', "000000000011000"),('1', "000000001010010"),('0', "000000000101010"),('1', "000000010001010"),('1', "000000000001010"),('1', "000000000111111"),('1', "000000000010001"),('1', "000000100111000")),
 ------------------------------- 
(('1', "000000000001000"),('1', "000000001001100"),('1', "000000000100111"),('1', "000000001001100"),('0', "000000000011001"),('1', "000000001001110"),('0', "000000000100010"),('0', "000000000010010"),('1', "000000000010001"),('0', "000000000111000"),('1', "000000000110101"),('0', "000000001000000"),('1', "000000010000110"),('1', "000000001100100"),('0', "000000000000101"),('1', "000000000010110"),('1', "000000001100111"),('1', "000000001111110"),('1', "000000011011100"),('0', "000000010010000"),('0', "000000001000100"),('1', "000000001010001"),('1', "000000001101001"),('1', "000000010111100"),('1', "000000010011101"),('0', "000000010101110"),('1', "000000000000110"),('1', "000000000110101"),('0', "000000011011110"),('1', "000000001111000"),('1', "000000000101110"),('0', "000000010010010"),('0', "000000001010101"),('1', "000000001100101"),('1', "000000000011011"),('0', "000000000110000"),('1', "000000000011111"),('1', "000000000110110"),('1', "000000001010101"),('0', "000000000100101"),('0', "000000000010001"),('0', "000000000111100"),('1', "000000001010111"),('0', "000000011000111"),('0', "000000000111011"),('0', "000000000111111"),('0', "000000001010100"),('0', "000000001000010"),('0', "000000011001000"),('0', "000000000000101"),('1', "000000000100110"),('0', "000000000000111"),('1', "000000000110000"),('0', "000000000010110"),('1', "000000000110110"),('1', "000000000101001"),('0', "000000000111000"),('1', "000000000110111"),('1', "000000001101110"),('1', "000000000111010"),('1', "000000001010111"),('1', "000000000101101"),('1', "000000100011111")),
 ------------------------------- 
(('1', "000000001011111"),('0', "000000000101100"),('0', "000000001100011"),('0', "000000000100011"),('1', "000000000001010"),('0', "000000000101001"),('1', "000000001000001"),('1', "000000000010101"),('1', "000000000011011"),('0', "000000000100110"),('1', "000000001010111"),('1', "000000010000101"),('0', "000000010110101"),('0', "000000001111001"),('1', "000000000110001"),('1', "000000000111010"),('1', "000000010011111"),('1', "000000000001000"),('1', "000000000111100"),('1', "000000001111110"),('0', "000000010010000"),('0', "000000001101000"),('0', "000000001100000"),('1', "000000001110101"),('1', "000000001110111"),('1', "000000011011100"),('1', "000000000100111"),('1', "000000011100101"),('1', "000000001001000"),('0', "000000000111110"),('1', "000000001011010"),('0', "000000000011010"),('1', "000000001100000"),('1', "000000001010100"),('0', "000000000010011"),('1', "000000001010010"),('1', "000000000000101"),('0', "000000000010011"),('0', "000000000001111"),('1', "000000010110011"),('1', "000000001100010"),('1', "000000001011011"),('1', "000000000010011"),('0', "000000011111001"),('0', "000000000000110"),('1', "000000001011000"),('0', "000000011001010"),('1', "000000001000010"),('1', "000000000101011"),('0', "000000001100000"),('1', "000000000100010"),('1', "000000001010010"),('0', "000000001001011"),('1', "000000000001101"),('0', "000000010111010"),('1', "000000000010010"),('1', "000000001110100"),('0', "000000000110010"),('0', "000000010010101"),('0', "000000000010010"),('0', "000000000110001"),('0', "000000001001110"),('0', "000000001101100")),
 ------------------------------- 
(('1', "000000001001010"),('1', "000000000010000"),('1', "000000001011111"),('1', "000000001100111"),('0', "000000000001001"),('0', "000000000000110"),('1', "000000000001101"),('1', "000000000101100"),('0', "000000001001101"),('0', "000000000101000"),('1', "000000000101100"),('1', "000000000010001"),('0', "000000000101000"),('0', "000000000100111"),('0', "000000000001110"),('0', "000000000101110"),('0', "000000000101000"),('1', "000000000011011"),('0', "000000000100110"),('0', "000000000111001"),('1', "000000001000000"),('1', "000000000001010"),('0', "000000000110000"),('0', "000000001000110"),('1', "000000000010010"),('0', "000000000100110"),('1', "000000000100000"),('0', "000000000001100"),('1', "000000100000101"),('1', "000000011100010"),('0', "000000000110111"),('0', "000000000001101"),('1', "000000001001010"),('0', "000000001000110"),('0', "000000000000110"),('0', "000000001100011"),('1', "000000010100000"),('0', "000000000101111"),('0', "000000000110000"),('0', "000000000111101"),('1', "000000000001101"),('0', "000000000010111"),('1', "000000001111011"),('1', "000000010100100"),('1', "000000000100111"),('0', "000000001000010"),('1', "000000000001010"),('0', "000000000011001"),('1', "000000001101100"),('0', "000000000000101"),('1', "000000000110101"),('1', "000000000100010"),('1', "000000000001011"),('0', "000000001000100"),('1', "000000000000101"),('1', "000000000001101"),('1', "000000001011011"),('0', "000000000010100"),('1', "000000000001110"),('0', "000000000101011"),('0', "000000000100111"),('1', "000000000001010"),('1', "000001000110010")),
 ------------------------------- 
(('1', "000000000100010"),('0', "000000000001010"),('1', "000000000100010"),('1', "000000000101010"),('0', "000000000000101"),('0', "000000000100101"),('1', "000000000100111"),('1', "000000000001000"),('0', "000000000110110"),('0', "000000001110011"),('0', "000000000111011"),('0', "000000001100010"),('0', "000000001000011"),('0', "000000000111100"),('0', "000000001000101"),('1', "000000000000111"),('0', "000000001001100"),('0', "000000001010101"),('0', "000000001000111"),('1', "000000000111110"),('0', "000000000000100"),('0', "000000000100101"),('0', "000000001110111"),('0', "000000000011111"),('1', "000000000111111"),('0', "000000001110010"),('1', "000000010111001"),('1', "000000000101000"),('1', "000000001001000"),('0', "000000000001000"),('1', "000000001000010"),('0', "000000000100111"),('1', "000000000111111"),('1', "000000000100010"),('1', "000000010101110"),('1', "000000001011101"),('1', "000000000110011"),('1', "000000000110100"),('0', "000000001111010"),('1', "000000011011000"),('1', "000000001110101"),('1', "000000000110110"),('1', "000000000000100"),('1', "000000000110001"),('1', "000000000001110"),('0', "000000000100000"),('1', "000000000010110"),('1', "000000000010111"),('1', "000000001010011"),('0', "000000001000110"),('0', "000000000100000"),('0', "000000001110011"),('0', "000000000110001"),('0', "000000001001100"),('0', "000000000110101"),('1', "000000000110111"),('1', "000000010001100"),('0', "000000001000101"),('0', "000000000110010"),('1', "000000000000001"),('0', "000000000111101"),('0', "000000000010001"),('0', "000000001110100")),
 ------------------------------- 
(('1', "000000001100010"),('1', "000000000000101"),('1', "000000011001000"),('0', "000000000000110"),('0', "000000000101110"),('0', "000000001000110"),('0', "000000001011101"),('1', "000000000011011"),('0', "000000000011110"),('0', "000000001010000"),('0', "000000000010100"),('0', "000000000100110"),('0', "000000010011011"),('0', "000000001000010"),('0', "000000000101100"),('1', "000000000000100"),('1', "000000000000111"),('0', "000000000101011"),('1', "000000000011001"),('1', "000000000101011"),('0', "000000000001111"),('0', "000000000110101"),('0', "000000000100000"),('1', "000000000010010"),('1', "000000000100100"),('1', "000000000001011"),('1', "000000000001010"),('0', "000000000000111"),('0', "000000000011000"),('0', "000000000010000"),('1', "000000000100001"),('0', "000000000100000"),('1', "000000000110100"),('0', "000000000001000"),('1', "000000000100001"),('0', "000000000100010"),('1', "000000000000011"),('1', "000000000011000"),('0', "000000000110001"),('1', "000000000011101"),('1', "000000000101011"),('1', "000000000010100"),('1', "000000001010000"),('1', "000000000100001"),('1', "000000010001011"),('0', "000000001000100"),('1', "000000001001000"),('0', "000000000000110"),('0', "000000000001111"),('0', "000000001100100"),('1', "000000001000011"),('1', "000000011100010"),('1', "000000000000110"),('1', "000000000101011"),('0', "000000000000010"),('1', "000000001001100"),('1', "000000010010111"),('0', "000000000001110"),('1', "000000000000101"),('1', "000000000101010"),('1', "000000001100001"),('1', "000000000000010"),('1', "000000111110000")),
 ------------------------------- 
(('1', "000000000101000"),('1', "000000001000111"),('0', "000000001101111"),('1', "000000000001011"),('1', "000000000000110"),('1', "000000000001100"),('0', "000000000011001"),('0', "000000001000011"),('0', "000000000000001"),('1', "000000010000000"),('0', "000000001110101"),('0', "000000010011101"),('1', "000000011001011"),('1', "000000010111010"),('1', "000000100110110"),('1', "000000110110001"),('0', "000000010111001"),('1', "000000010000011"),('0', "000000000000110"),('0', "000000000010001"),('0', "000000000000101"),('0', "000000000110011"),('0', "000000001000011"),('1', "000000010011011"),('0', "000000000000101"),('1', "000000000000011"),('0', "000000000100000"),('0', "000000000001100"),('0', "000000000010000"),('0', "000000000000001"),('0', "000000000101000"),('1', "000000010011101"),('0', "000000001010010"),('1', "000000000001100"),('0', "000000000000111"),('1', "000000001101100"),('1', "000000000101111"),('1', "000000001000111"),('0', "000000000010111"),('1', "000000000001010"),('1', "000000000000110"),('0', "000000001111111"),('0', "000000000110100"),('0', "000000001100110"),('1', "000000000100101"),('0', "000000001111100"),('0', "000000000010001"),('1', "000000000101001"),('1', "000000001001010"),('1', "000000000010110"),('1', "000000000010010"),('0', "000000011001010"),('0', "000000001011011"),('1', "000000000010110"),('0', "000000001000011"),('1', "000000000010100"),('1', "000000000010001"),('1', "000000010010000"),('1', "000000000001001"),('1', "000000001100101"),('0', "000000000011000"),('1', "000000000000100"),('1', "000000100000100")),
 ------------------------------- 
(('1', "000000001000011"),('0', "000000001000111"),('1', "000000000110001"),('0', "000000000000000"),('0', "000000001001010"),('0', "000000000010000"),('1', "000000000001100"),('1', "000000000001010"),('1', "000000000110000"),('0', "000000000010010"),('1', "000000000100011"),('1', "000000000011101"),('1', "000000000011111"),('1', "000000000010001"),('0', "000000001010011"),('0', "000000001111101"),('1', "000000010110111"),('1', "000000001000100"),('1', "000000000111011"),('0', "000000010101110"),('1', "000000000101000"),('1', "000000001101101"),('0', "000000000000111"),('0', "000000010011010"),('1', "000000010110001"),('0', "000000001001100"),('0', "000000000111011"),('1', "000000000010010"),('0', "000000000000101"),('0', "000000000100011"),('1', "000000001010110"),('1', "000000000101100"),('0', "000000000011110"),('0', "000000010100000"),('1', "000000000101010"),('0', "000000000001001"),('1', "000000001111011"),('1', "000000001011011"),('1', "000000000100011"),('0', "000000010010100"),('1', "000000000010000"),('1', "000000010000110"),('1', "000000000000011"),('1', "000000000011100"),('1', "000000000000010"),('0', "000000000011000"),('0', "000000010101011"),('0', "000000001010110"),('0', "000000000101111"),('1', "000000000100110"),('0', "000000000100100"),('0', "000000000010001"),('1', "000000000000001"),('1', "000000000011010"),('1', "000000000011111"),('0', "000000001000110"),('0', "000000001101000"),('1', "000000001000001"),('0', "000000000000111"),('0', "000000010011100"),('0', "000000000001111"),('0', "000000000100110"),('0', "000000000101011")),
 ------------------------------- 
(('1', "000000001011011"),('1', "000000011100001"),('1', "000000000100110"),('0', "000000000000101"),('0', "000000000011011"),('1', "000000001101010"),('1', "000000000000011"),('1', "000000000011110"),('1', "000000000011010"),('0', "000000000001111"),('0', "000000000000001"),('1', "000000000001000"),('1', "000000000011100"),('1', "000000000001001"),('1', "000000000001011"),('1', "000000000101010"),('1', "000000001011011"),('1', "000000000001011"),('0', "000000000010011"),('1', "000000000001100"),('0', "000000010000100"),('0', "000000000011111"),('1', "000000000111110"),('0', "000000000101110"),('1', "000000000000001"),('1', "000000001100010"),('0', "000000000100000"),('1', "000000000011010"),('0', "000000000111000"),('0', "000000001010101"),('0', "000000000100110"),('0', "000000000001010"),('1', "000000001000010"),('1', "000000000000101"),('0', "000000001010111"),('0', "000000001101011"),('0', "000000000101110"),('0', "000000000011010"),('1', "000000001101111"),('1', "000000001000001"),('0', "000000010000001"),('0', "000000001110000"),('1', "000000000100001"),('0', "000000000101100"),('1', "000000001011011"),('1', "000000000110010"),('0', "000000000100011"),('0', "000000000001111"),('1', "000000000100110"),('1', "000000000010101"),('1', "000000001001000"),('1', "000000011100110"),('1', "000000000010110"),('1', "000000001011111"),('1', "000000000011110"),('0', "000000000000000"),('1', "000000001101000"),('0', "000000000010111"),('1', "000000000000111"),('1', "000000000100001"),('1', "000000000011011"),('0', "000000000100111"),('1', "000001000001000")),
 ------------------------------- 
(('1', "000000000110100"),('0', "000000000100110"),('0', "000000000011011"),('0', "000000001010010"),('1', "000000000100011"),('0', "000000001101010"),('1', "000000001000011"),('1', "000000000101101"),('1', "000000000101001"),('0', "000000000111001"),('0', "000000001110011"),('1', "000000000010001"),('0', "000000010010001"),('0', "000000000110011"),('0', "000000001000111"),('0', "000000000111011"),('0', "000000001101100"),('0', "000000011110111"),('0', "000000001100100"),('1', "000000000101110"),('1', "000000000001000"),('1', "000000000011110"),('1', "000000000100000"),('1', "000000011100111"),('1', "000000000101101"),('0', "000000000100011"),('1', "000000001111110"),('1', "000000000000011"),('1', "000000000011111"),('0', "000000000110111"),('1', "000000011011100"),('1', "000000001010100"),('0', "000000000001111"),('1', "000000000001000"),('0', "000000000011100"),('1', "000000000101011"),('1', "000000000010101"),('0', "000000000100000"),('0', "000000000001100"),('1', "000000000100110"),('1', "000000001110101"),('1', "000000100110000"),('0', "000000000101011"),('1', "000000001001000"),('1', "000000000000011"),('0', "000000001000010"),('0', "000000010000110"),('0', "000000010011000"),('0', "000000001100100"),('0', "000000001000100"),('0', "000000001100001"),('0', "000000010111110"),('0', "000000001100111"),('0', "000000000010010"),('0', "000000001100000"),('0', "000000001000101"),('0', "000000000100101"),('0', "000000001010110"),('1', "000000000010101"),('0', "000000001011100"),('1', "000000000101110"),('0', "000000000001001"),('0', "000000010100111")),
 ------------------------------- 
(('1', "000000000101110"),('0', "000000001001100"),('1', "000000001001111"),('0', "000000000100111"),('0', "000000000000010"),('1', "000000000101000"),('1', "000000001100011"),('1', "000000010011010"),('1', "000000010100111"),('1', "000000000010101"),('1', "000000000000001"),('1', "000000000000100"),('0', "000000001101111"),('1', "000000010101000"),('1', "000000011010000"),('1', "000000001011101"),('1', "000000000110101"),('0', "000000000000111"),('0', "000000010100111"),('1', "000000000001111"),('1', "000000010101101"),('1', "000000001101111"),('1', "000000000101000"),('1', "000000000001011"),('0', "000000000010101"),('0', "000000001011011"),('1', "000000010000100"),('0', "000000000010001"),('0', "000000000001001"),('0', "000000000111010"),('0', "000000000011000"),('0', "000000000010111"),('0', "000000000000001"),('0', "000000000101000"),('1', "000000001000000"),('1', "000000010000001"),('1', "000000001000100"),('0', "000000001011011"),('0', "000000001111100"),('1', "000000001100011"),('0', "000000000111011"),('1', "000000010001111"),('0', "000000100000101"),('0', "000000001101100"),('0', "000000000100011"),('0', "000000001101111"),('0', "000000001010000"),('0', "000000010001011"),('0', "000000000001100"),('1', "000000001001001"),('0', "000000010111101"),('0', "000000001000110"),('0', "000000001111111"),('0', "000000000000110"),('0', "000000011011101"),('0', "000000000010100"),('0', "000000000100110"),('1', "000000001101001"),('1', "000000000100111"),('1', "000000000000001"),('1', "000000000101111"),('1', "000000001001000"),('1', "000000010010000")),
 ------------------------------- 
(('0', "000000000000101"),('1', "000000000000010"),('0', "000000000101110"),('1', "000000001111000"),('1', "000000000111000"),('1', "000000010100100"),('1', "000000000110101"),('1', "000000000001100"),('0', "000000001011110"),('0', "000000000110001"),('0', "000000010100000"),('1', "000000010010011"),('0', "000000001111011"),('1', "000000000100001"),('0', "000000000101011"),('1', "000000010010001"),('0', "000000010010001"),('0', "000000000100000"),('0', "000000000110010"),('1', "000000010110111"),('0', "000000000111101"),('0', "000000010110111"),('0', "000000001001100"),('1', "000000011010001"),('0', "000000001100001"),('1', "000000001100000"),('0', "000000001111111"),('0', "000000110101010"),('1', "000000000100001"),('1', "000000000000010"),('1', "000000100100111"),('0', "000000000011011"),('0', "000000001100000"),('0', "000000011010000"),('1', "000000011010011"),('0', "000000000110101"),('0', "000000000100001"),('1', "000000000100010"),('0', "000000001011111"),('0', "000000100010111"),('1', "000000010001100"),('0', "000000010011111"),('1', "000000000100110"),('0', "000000000111001"),('1', "000000001111100"),('0', "000000001110101"),('1', "000000001111101"),('0', "000000011110011"),('1', "000000001000001"),('0', "000000011001110"),('1', "000000011111001"),('0', "000000011000001"),('0', "000000001011101"),('0', "000000001000011"),('1', "000000001000001"),('0', "000000000000100"),('0', "000000001111100"),('0', "000000100010010"),('1', "000000010010011"),('0', "000000000011000"),('0', "000000001000001"),('1', "000000001010100"),('1', "000000000010010")),
 ------------------------------- 
(('0', "000000010000000"),('1', "000000000111101"),('0', "000000000100111"),('1', "000000001110111"),('0', "000000000110110"),('0', "000000000011100"),('1', "000000000100001"),('0', "000000000111110"),('0', "000000000000100"),('0', "000000000000001"),('1', "000000000010000"),('0', "000000000011011"),('1', "000000000001110"),('0', "000000000100000"),('0', "000000000001000"),('0', "000000001010100"),('0', "000000001101001"),('0', "000000000000011"),('0', "000000001010101"),('0', "000000001000101"),('1', "000000000000111"),('0', "000000000000010"),('0', "000000000100011"),('0', "000000000001100"),('0', "000000001101111"),('1', "000000001110111"),('1', "000000010001111"),('0', "000000001010001"),('0', "000000000111101"),('1', "000000001000000"),('1', "000000000011110"),('1', "000000010000001"),('1', "000000010110000"),('1', "000000001000100"),('1', "000000000111010"),('1', "000000001000011"),('1', "000000000010110"),('0', "000000000001010"),('1', "000000011100100"),('0', "000000000010001"),('1', "000000001100000"),('1', "000000001011110"),('0', "000000001111110"),('1', "000000001100101"),('1', "000000001010001"),('1', "000000001010100"),('0', "000000000000101"),('0', "000000000000110"),('0', "000000000100011"),('1', "000000001000001"),('0', "000000001010111"),('0', "000000010000101"),('0', "000000001000010"),('0', "000000000010000"),('1', "000000000111110"),('0', "000000001000101"),('1', "000000001000110"),('1', "000000001001010"),('1', "000000001100000"),('0', "000000000010001"),('0', "000000000001000"),('1', "000000001110000"),('1', "000000011010000")),
 ------------------------------- 
(('0', "000000101010101"),('1', "000000000010001"),('0', "000000000111000"),('1', "000000011111100"),('1', "000000000100000"),('0', "000000000100011"),('1', "000000000011111"),('0', "000000010000000"),('0', "000000001101000"),('1', "000000000111000"),('1', "000000010001000"),('1', "000000001000001"),('0', "000000000110011"),('0', "000000010100101"),('1', "000000000111011"),('0', "000000010001110"),('0', "000000000000100"),('1', "000000000010110"),('0', "000000001100010"),('1', "000000010000100"),('0', "000000010000000"),('0', "000000010110001"),('1', "000000001011100"),('0', "000000001001001"),('0', "000000000011011"),('1', "000000001111101"),('0', "000000001001101"),('0', "000000010011100"),('1', "000000000000011"),('0', "000000001110001"),('0', "000000011101100"),('1', "000000010011110"),('1', "000000000010011"),('0', "000000001100110"),('0', "000000000111101"),('1', "000000000100010"),('0', "000000000100011"),('0', "000000000001110"),('0', "000000001100010"),('0', "000000001110110"),('1', "000000000010010"),('0', "000000001010111"),('0', "000000000000100"),('1', "000000100000011"),('1', "000000010001010"),('0', "000000000011010"),('1', "000000010010101"),('1', "000000000100001"),('1', "000000010011111"),('1', "000000001111011"),('1', "000000000101100"),('0', "000000000000100"),('0', "000000000110111"),('1', "000000000100101"),('1', "000000001011000"),('0', "000000001100101"),('1', "000000000101111"),('1', "000000001011010"),('1', "000000001011000"),('0', "000000000010000"),('1', "000000000000010"),('1', "000000001011010"),('0', "000000100010110")),
 ------------------------------- 
(('0', "000000000111001"),('0', "000000000101001"),('0', "000000000001010"),('0', "000000001010101"),('1', "000000001001011"),('0', "000000001010001"),('0', "000000000110010"),('0', "000000000000101"),('1', "000000000000010"),('1', "000000000010101"),('0', "000000010111101"),('1', "000000000110111"),('0', "000000010101111"),('1', "000000001000101"),('0', "000000001000110"),('0', "000000000011101"),('1', "000000000011000"),('0', "000000000111000"),('0', "000000000011001"),('1', "000000001000100"),('1', "000000000001010"),('1', "000000001001000"),('1', "000000000100010"),('1', "000000010110010"),('1', "000000010000101"),('1', "000000000110101"),('1', "000000000001111"),('0', "000000000000110"),('1', "000000001011110"),('1', "000000000110101"),('1', "000000001001111"),('0', "000000001101100"),('1', "000000001001100"),('1', "000000000100100"),('1', "000000001010011"),('0', "000000000110001"),('1', "000000000010001"),('0', "000000001101011"),('1', "000000001100010"),('0', "000000001001101"),('1', "000000000100110"),('1', "000000000010010"),('1', "000000001011100"),('1', "000000101010101"),('0', "000000001000001"),('0', "000000000100110"),('1', "000000001111111"),('0', "000000001001001"),('0', "000000000100110"),('1', "000000000101111"),('0', "000000010000110"),('0', "000000000110111"),('0', "000000000011110"),('1', "000000000010100"),('1', "000000000000101"),('1', "000000000010011"),('0', "000000001001010"),('1', "000000000011011"),('0', "000000000011010"),('1', "000000000110000"),('1', "000000000110010"),('1', "000000000011100"),('1', "000000010100100")),
 ------------------------------- 
(('0', "000000000011110"),('1', "000000000100010"),('1', "000000000000011"),('0', "000000001101101"),('0', "000000000101010"),('0', "000000000100111"),('0', "000000000011010"),('1', "000000000001110"),('0', "000000000001101"),('1', "000000001010010"),('0', "000000000010111"),('0', "000000001000101"),('1', "000000000100111"),('0', "000000000011111"),('0', "000000000001000"),('1', "000000000100000"),('1', "000000011011110"),('1', "000000011111010"),('1', "000000011111111"),('1', "000000000001011"),('1', "000000000100100"),('0', "000000000010011"),('0', "000000001110000"),('0', "000000000011010"),('0', "000000000111000"),('0', "000000001100100"),('0', "000000000100010"),('1', "000000000101010"),('1', "000000001101000"),('1', "000000010000011"),('1', "000000000010000"),('0', "000000000000001"),('0', "000000000100010"),('0', "000000001110010"),('1', "000000000101011"),('0', "000000001010011"),('0', "000000000010100"),('1', "000000000011011"),('1', "000000001000011"),('0', "000000001010110"),('1', "000000000101111"),('0', "000000001010100"),('1', "000000000011000"),('0', "000000001001011"),('0', "000000000100110"),('0', "000000001000100"),('1', "000000000101011"),('1', "000000000000111"),('1', "000000000100010"),('0', "000000000101110"),('1', "000000000111111"),('1', "000000000011101"),('1', "000000000001111"),('0', "000000010000010"),('0', "000000000001010"),('1', "000000000110001"),('1', "000000000001011"),('0', "000000000110000"),('0', "000000001001001"),('0', "000000000111111"),('0', "000000001000101"),('0', "000000001101111"),('1', "000000000011000")),
 ------------------------------- 
(('1', "000000000001011"),('0', "000000000000001"),('0', "000000000010101"),('0', "000000001011010"),('0', "000000000001101"),('0', "000000000011000"),('1', "000000000010110"),('0', "000000000000111"),('1', "000000000001111"),('1', "000000000010000"),('0', "000000000100111"),('0', "000000001011011"),('0', "000000000100100"),('0', "000000000101001"),('0', "000000000010010"),('0', "000000000101100"),('1', "000000010111101"),('1', "000000001111101"),('0', "000000000011111"),('0', "000000010010001"),('1', "000000000000100"),('1', "000000000111001"),('0', "000000000001000"),('0', "000000000011111"),('1', "000000010001010"),('0', "000000000101010"),('0', "000000010111111"),('1', "000000001011010"),('0', "000000000100000"),('1', "000000000101011"),('1', "000000000100100"),('1', "000000000011101"),('0', "000000001001010"),('0', "000000001001111"),('1', "000000000001010"),('1', "000000000111001"),('1', "000000000000110"),('1', "000000011101111"),('1', "000000011101000"),('0', "000000001010000"),('1', "000000000100100"),('1', "000000000111000"),('0', "000000000001011"),('1', "000000000001011"),('1', "000000000010110"),('1', "000000010101010"),('1', "000000010111110"),('0', "000000000000111"),('1', "000000000111010"),('1', "000000000111001"),('0', "000000001001001"),('1', "000000000110100"),('1', "000000000011110"),('0', "000000000001001"),('1', "000000000101101"),('0', "000000000011100"),('1', "000000000010110"),('1', "000000000010100"),('0', "000000001000110"),('1', "000000000000101"),('0', "000000000111111"),('1', "000000000000110"),('0', "000000000001011")),
 ------------------------------- 
(('1', "000000001000101"),('0', "000000000100100"),('0', "000000010000100"),('1', "000000000000101"),('1', "000000001000101"),('1', "000000001100101"),('1', "000000001111001"),('1', "000000010011101"),('1', "000000000001001"),('1', "000000000000010"),('0', "000000001110000"),('0', "000000000000111"),('0', "000000000001101"),('0', "000000000011011"),('1', "000000000010011"),('0', "000000010000111"),('1', "000000001011111"),('0', "000000001000101"),('0', "000000000110010"),('0', "000000010110011"),('0', "000000001001100"),('0', "000000000100111"),('0', "000000000010100"),('1', "000000000111110"),('1', "000000000110011"),('1', "000000000001011"),('1', "000000000111101"),('1', "000000000100110"),('1', "000000000100110"),('1', "000000001111000"),('0', "000000000011100"),('1', "000000000010000"),('1', "000000000011101"),('1', "000000001011101"),('1', "000000000100010"),('0', "000000000100111"),('1', "000000001010000"),('1', "000000000111001"),('1', "000000000010100"),('1', "000000000100110"),('0', "000000001011011"),('0', "000000001111101"),('0', "000000000011101"),('0', "000000001110111"),('0', "000000000101101"),('0', "000000000100100"),('1', "000000000011001"),('1', "000000000011011"),('1', "000000000111110"),('1', "000000001000001"),('0', "000000000010010"),('0', "000000001000101"),('1', "000000000011101"),('0', "000000000001001"),('1', "000000001110000"),('0', "000000000101001"),('1', "000000000110011"),('1', "000000001100010"),('1', "000000001000001"),('0', "000000000010000"),('0', "000000001001100"),('1', "000000000110110"),('1', "000000100010000"))
 ------------------------------- 
);	
begin
	process(clk) 
	begin -- process
		if clk'event and clk = '1' then
			if (en = '1') then
				for i in 0 to address_size-1 LOOP
					ROM_data(i) <= rom(i)(address);
				end LOOP;
			end if;
		end if;
	end process;
end weight_L1;

architecture weight_L2 of ROM is

	type rom_type is array (0 to address_size-1) of fixed_point_array (0 to entry_length-1);
	signal rom : rom_type:=(
(('0', "000000000000000"),('0', "000000000000001"),('1', "000000000000010"),('1', "000000000000011"),('0', "000000000000000"),('1', "000000000001010"),('0', "000000000000011"),('1', "000000000000001"),('1', "000000000000010"),('0', "000000000000001"),('1', "000000000000111"),('1', "000000000000100"),('1', "000000000000001"),('0', "000000000000000"),('1', "000000000000001"),('1', "000000000000001"),('0', "000000000000000"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000011")),
----------------------------
(('0', "000000000000100"),('1', "000000000000111"),('0', "000000000000000"),('0', "000000000000100"),('0', "000000000000011"),('0', "000000000000101"),('1', "000000000001000"),('1', "000000000000101"),('0', "000000000000010"),('0', "000000000000001"),('0', "000000000000001"),('0', "000000000000010"),('0', "000000000000000"),('0', "000000000000010"),('0', "000000000000100"),('0', "000000000000010"),('0', "000000000000000"),('1', "000000000000101"),('0', "000000000000011"),('1', "000000000000100")),
----------------------------
(('1', "000000000000001"),('1', "000000000000010"),('0', "000000000000011"),('0', "000000000000011"),('0', "000000000000010"),('1', "000000000000111"),('1', "000000000000011"),('0', "000000000000000"),('0', "000000000000001"),('0', "000000000000000"),('1', "000000000000101"),('0', "000000000000010"),('1', "000000000000100"),('1', "000000000000010"),('1', "000000000000001"),('0', "000000000000010"),('0', "000000000000011"),('0', "000000000000010"),('1', "000000000000100"),('0', "000000000000010")),
----------------------------
(('1', "000000000000010"),('0', "000000000000000"),('1', "000000000000011"),('0', "000000000000001"),('1', "000000000000001"),('1', "000000000000100"),('1', "000000000000011"),('0', "000000000000001"),('1', "000000000000100"),('1', "000000000000100"),('1', "000000000000101"),('1', "000000000000001"),('0', "000000000000010"),('0', "000000000000001"),('0', "000000000000010"),('0', "000000000000000"),('1', "000000000000010"),('0', "000000000000001"),('0', "000000000000100"),('0', "000000000000000")),
----------------------------
(('1', "000000000000001"),('1', "000000000000001"),('0', "000000000000011"),('1', "000000000000001"),('1', "000000000000011"),('0', "000000000000000"),('1', "000000000001000"),('1', "000000000001100"),('1', "000000000000100"),('1', "000000000000011"),('0', "000000000000010"),('1', "000000000001000"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000001"),('1', "000000000000110"),('1', "000000000000001"),('1', "000000000001001")),
----------------------------
(('0', "000000000000100"),('0', "000000000000000"),('1', "000000000000100"),('0', "000000000000000"),('1', "000000000000001"),('0', "000000000001000"),('1', "000000000000101"),('0', "000000000000001"),('0', "000000000000010"),('1', "000000000000110"),('1', "000000000001000"),('0', "000000000000010"),('1', "000000000000011"),('1', "000000000000010"),('1', "000000000000001"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000010"),('0', "000000000000000"),('0', "000000000000110")),
----------------------------
(('1', "000000000000001"),('1', "000000000000001"),('1', "000000000000100"),('0', "000000000000000"),('0', "000000000000000"),('0', "000000000000010"),('1', "000000000000010"),('1', "000000000000001"),('0', "000000000000001"),('0', "000000000000000"),('1', "000000000000001"),('1', "000000000000100"),('0', "000000000000100"),('0', "000000000000000"),('0', "000000000000000"),('1', "000000000000010"),('1', "000000000000001"),('1', "000000000000010"),('1', "000000000000011"),('1', "000000000000100")),
----------------------------
(('1', "000000000000011"),('1', "000000000000100"),('0', "000000000000010"),('1', "000000000000001"),('0', "000000000000001"),('0', "000000000000100"),('1', "000000000000011"),('0', "000000000000011"),('0', "000000000000010"),('1', "000000000000001"),('0', "000000000000101"),('1', "000000000000010"),('1', "000000000000011"),('0', "000000000000001"),('0', "000000000000111"),('1', "000000000000011"),('0', "000000000000010"),('0', "000000000000010"),('1', "000000000000001"),('1', "000000000000010")),
----------------------------
(('1', "000000000001001"),('1', "000000000000110"),('1', "000000000000010"),('1', "000000000000110"),('1', "000000000000111"),('1', "000000000000010"),('0', "000000000000011"),('1', "000000000000011"),('0', "000000000000001"),('0', "000000000000011"),('1', "000000000001001"),('1', "000000000000010"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000101"),('1', "000000000000010"),('0', "000000000000010"),('1', "000000000000011"),('1', "000000000000010"),('1', "000000000000011")),
----------------------------
(('1', "000000000000110"),('0', "000000000000010"),('1', "000000000000011"),('1', "000000000000010"),('1', "000000000000001"),('0', "000000000000001"),('1', "000000000000111"),('0', "000000000001000"),('0', "000000000000001"),('1', "000000000000101"),('1', "000000000000011"),('1', "000000000000001"),('1', "000000000000100"),('1', "000000000000010"),('1', "000000000000111"),('1', "000000000000001"),('1', "000000000001001"),('1', "000000000000110"),('0', "000000000000001"),('1', "000000000000010"))
);	
begin
	process(clk) 
	begin -- process
		if clk'event and clk = '1' then
			if (en = '1') then
				for i in 0 to address_size-1 LOOP
					ROM_data(i) <= rom(i)(address);
				end LOOP;
			end if;
		end if;
	end process;
end weight_L2;

architecture weight_test1 of ROM is
	type rom_type is array (0 to address_size-1) of fixed_point_array (0 to entry_length-1);
	signal rom : rom_type:=(
	
		(('0', "000000000000000"),('0', "000000001000000"),('0', "000000010000000"),('0', "000000000000000")), ----- 0, 1, 2, 0
		------------------------------- 
		(('0', "000000001000000"),('0', "000000000000000"),('0', "000000000000000"),('0', "000000011000000")) ----- 1, 0, 0, 3
		------------------------------- 
	);
begin
	process(clk) 
	begin -- process
		if clk'event and clk = '1' then
			if (en = '1') then
				for i in 0 to address_size-1 LOOP
					ROM_data(i) <= rom(i)(address);
				end LOOP;
			end if;
		end if;
	end process;
end weight_test1;

architecture weight_test2 of ROM is
	type rom_type is array (0 to address_size-1) of fixed_point_array (0 to entry_length-1);
	signal rom : rom_type:=(
	
		(('0', "000000000000000"),('0', "000000001000000")), ----- 0, 1
		------------------------------- 
		(('0', "000000001000000"),('0', "000000000000000")) ----- 1, 0
		------------------------------- 
	);
begin
	process(clk) 
	begin -- process
		if clk'event and clk = '1' then
			if (en = '1') then
				for i in 0 to address_size-1 LOOP
					ROM_data(i) <= rom(i)(address);
				end LOOP;
			end if;
		end if;
	end process;
end weight_test2;
